module mux4way16(
    input[15:0] a,
    input[15:0] b,
    input[15:0] c,
    input[15:0] d,
    input[1:0] sel,
    output[15:0] out
);
endmodule
