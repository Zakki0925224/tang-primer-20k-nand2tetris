`default_nettype none

module not16(
    input wire[15:0] in,
    output wire[15:0] out
);
    _not not_gate_0(
        .in(in[0]),
        .out(out[0])
    );
    _not not_gate_1(
        .in(in[1]),
        .out(out[1])
    );
    _not not_gate_2(
        .in(in[2]),
        .out(out[2])
    );
    _not not_gate_3(
        .in(in[3]),
        .out(out[3])
    );
    _not not_gate_4(
        .in(in[4]),
        .out(out[4])
    );
    _not not_gate_5(
        .in(in[5]),
        .out(out[5])
    );
    _not not_gate_6(
        .in(in[6]),
        .out(out[6])
    );
    _not not_gate_7(
        .in(in[7]),
        .out(out[7])
    );
    _not not_gate_8(
        .in(in[8]),
        .out(out[8])
    );
    _not not_gate_9(
        .in(in[9]),
        .out(out[9])
    );
    _not not_gate_10(
        .in(in[10]),
        .out(out[10])
    );
    _not not_gate_11(
        .in(in[11]),
        .out(out[11])
    );
    _not not_gate_12(
        .in(in[12]),
        .out(out[12])
    );
    _not not_gate_13(
        .in(in[13]),
        .out(out[13])
    );
    _not not_gate_14(
        .in(in[14]),
        .out(out[14])
    );
    _not not_gate_15(
        .in(in[15]),
        .out(out[15])
    );
endmodule

`default_nettype wire
